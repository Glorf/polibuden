library verilog;
use verilog.vl_types.all;
entity Cwiczenie5_5_vlg_vec_tst is
end Cwiczenie5_5_vlg_vec_tst;
