library verilog;
use verilog.vl_types.all;
entity Cwiczenie5_1_vlg_sample_tst is
    port(
        iSW             : in     vl_logic_vector(0 to 3);
        sampler_tx      : out    vl_logic
    );
end Cwiczenie5_1_vlg_sample_tst;
