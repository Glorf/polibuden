library verilog;
use verilog.vl_types.all;
entity Cwiczenie3_4_vlg_check_tst is
    port(
        oLEDG           : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end Cwiczenie3_4_vlg_check_tst;
