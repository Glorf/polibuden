library verilog;
use verilog.vl_types.all;
entity Cwiczenie2_1_vlg_check_tst is
    port(
        oLEDG           : in     vl_logic_vector(2 downto 0);
        sampler_rx      : in     vl_logic
    );
end Cwiczenie2_1_vlg_check_tst;
