library verilog;
use verilog.vl_types.all;
entity Cwiczenie5_2_vlg_vec_tst is
end Cwiczenie5_2_vlg_vec_tst;
