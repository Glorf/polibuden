library verilog;
use verilog.vl_types.all;
entity Cwiczenie5_1_vlg_check_tst is
    port(
        oLEDG           : in     vl_logic_vector(0 to 1);
        sampler_rx      : in     vl_logic
    );
end Cwiczenie5_1_vlg_check_tst;
