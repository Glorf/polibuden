library verilog;
use verilog.vl_types.all;
entity Cwiczenie4_vlg_vec_tst is
end Cwiczenie4_vlg_vec_tst;
