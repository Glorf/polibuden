library verilog;
use verilog.vl_types.all;
entity Cwiczenie5_2_vlg_check_tst is
    port(
        sout            : in     vl_logic;
        sum             : in     vl_logic_vector(0 to 7);
        sampler_rx      : in     vl_logic
    );
end Cwiczenie5_2_vlg_check_tst;
