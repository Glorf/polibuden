library ieee;
use ieee.std_logic_1164.all;

entity char7seg is
	port(
		C: in std_logic_vector(2 downto 0);
		Display: out std_logic_vector(2 downto 0));
end char7seg;

architecture strukturalna of char7seg is
begin
--UZUPEŁNIĆ!
end strukturalna;