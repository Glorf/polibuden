library verilog;
use verilog.vl_types.all;
entity Cwiczenie5_1 is
    port(
        iSW             : in     vl_logic_vector(0 to 3);
        oLEDG           : out    vl_logic_vector(0 to 1)
    );
end Cwiczenie5_1;
