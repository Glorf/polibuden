library ieee;
use ieee.std_logic_1164.all;

entity Cwiczenie7 is
	Port(
		KEY: in std_logic_vector(0 to 1);
		LEDR: out std_logic_vector(0 to 0);
		SRAM_ADDR: in std_logic_vector(0 to 17);
		SRAM_DQ: 
	);
end Cwiczenie7;

architecture pamiec of Cwiczenie7 is
