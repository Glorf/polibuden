library verilog;
use verilog.vl_types.all;
entity Cwiczenie3_2_vlg_sample_tst is
    port(
        iSW             : in     vl_logic_vector(1 downto 0);
        sampler_tx      : out    vl_logic
    );
end Cwiczenie3_2_vlg_sample_tst;
