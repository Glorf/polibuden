library verilog;
use verilog.vl_types.all;
entity Cwiczenie3_2_vlg_vec_tst is
end Cwiczenie3_2_vlg_vec_tst;
