library verilog;
use verilog.vl_types.all;
entity Cwiczenie5_5_vlg_check_tst is
    port(
        w               : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end Cwiczenie5_5_vlg_check_tst;
