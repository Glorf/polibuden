library verilog;
use verilog.vl_types.all;
entity Cwiczenie3_4_vlg_sample_tst is
    port(
        iSW             : in     vl_logic_vector(2 downto 0);
        sampler_tx      : out    vl_logic
    );
end Cwiczenie3_4_vlg_sample_tst;
