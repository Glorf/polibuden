library verilog;
use verilog.vl_types.all;
entity Cwiczenie2_1_vlg_vec_tst is
end Cwiczenie2_1_vlg_vec_tst;
