library verilog;
use verilog.vl_types.all;
entity Cwiczenie5_3_vlg_check_tst is
    port(
        out0            : in     vl_logic_vector(0 to 7);
        overf           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Cwiczenie5_3_vlg_check_tst;
