library ieee;
use ieee.std_logic_1164.all;

entity mux3bit8to1 is
	port (
		S,U0,U1,U2,U3,U4,U5,U6,U7: in std_logic_vector(2 downto 0);
		M: out std_logic_vector(2 downto 0));
end mux3bit8to1;


architecture strukturalna of mux3bit8to1 is
begin
--UZUPEŁNIĆ
end strukturalna;