library verilog;
use verilog.vl_types.all;
entity Cwiczenie5_3_vlg_vec_tst is
end Cwiczenie5_3_vlg_vec_tst;
