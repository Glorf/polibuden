library verilog;
use verilog.vl_types.all;
entity Cwiczenie2_3_vlg_check_tst is
    port(
        oLEDG           : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end Cwiczenie2_3_vlg_check_tst;
