library verilog;
use verilog.vl_types.all;
entity Cwiczenie2_3_vlg_vec_tst is
end Cwiczenie2_3_vlg_vec_tst;
