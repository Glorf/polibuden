library verilog;
use verilog.vl_types.all;
entity Cwiczenie2_2_vlg_sample_tst is
    port(
        iSW             : in     vl_logic_vector(2 downto 0);
        sampler_tx      : out    vl_logic
    );
end Cwiczenie2_2_vlg_sample_tst;
